module tb_top;

    initial begin
        $display("Hello");
    end

endmodule
